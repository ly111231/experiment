module our;
	initial begin ("Hello World");
	$finish;
	end
		 
endmodule
